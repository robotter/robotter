-----------------------------------------------------------------------------
-- Title      : Threshold bloc
-- Project    : Carte camera 2009
-----------------------------------------------------------------------------
-- File       : threshold.vhdl
-- Author     : BLANCHARD Remy <remyb718 at gmail dot com>
-- Company    : Rob'Otter
-- Last update: 16/11/2008
-- Platform   : Spartan 3
-----------------------------------------------------------------------------
-- Description: Determine if the input are in or outside the wanted values
--              This bloc uses a block RAM per entry and a "AND" door: the 
--              value must within range for all inputs
-----------------------------------------------------------------------------
-- This program is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 2, or (at your option)
-- any later version.
-- 
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License
-- along with this program; if not, write to the Free Software
-----------------------------------------------------------------------------
-- HISTORY :
-- +------------------------------------------------------------------------+
-- | Ver. | Date     | Aut. | Commentaire                                   |
-- +------------------------------------------------------------------------+
-- | 1.00 | 16/11/08 | RBL  | Creation                                      |
-- +------------------------------------------------------------------------+
-- | 1.05 | 18/01/09 | RBL  | Modification of the H's output size           |
-- +------------------------------------------------------------------------+
-- |      |          |      |                                               |
-- +------------------------------------------------------------------------+
-- |      |          |      |                                               |
-- +------------------------------------------------------------------------+

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VComponents.all;

-----------------------------------------------------------------------
entity threshold is
-----------------------------------------------------------------------
    port (
        clk_i          : in  std_ulogic;
        -- input to be tested
        Y_i            : in  std_logic_vector(7 downto 0);
        H_i            : in  std_logic_vector(7 downto 0);

        -- threshold modifier (modify bloc RAM inside)
        valid_i        : in  std_ulogic; -- write RAM if active
		  value_i        : in  std_logic_vector(15 downto 0);
		  -- for adress_i: MSB=1 modify Y Look-Up Table else H LUT
        adress_i       : in  std_logic_vector(9 downto 0); 

        -- vector of all threshold result
        result_o       : out std_logic_vector(15 downto 0) --latched
    );
end threshold;

-----------------------------------------------------------------------
architecture threshold_1 of threshold is
-----------------------------------------------------------------------

-- declaration

    -- Y memory signals
    signal Y_thres_s    : std_logic_vector(15 downto 0);
    signal Y_ADDR_A_s   : std_logic_vector(9 downto 0);
    signal Y_ADDR_B_s   : std_logic_vector(9 downto 0);
    signal Y_enable_B_s : std_ulogic;

    signal H_thres_s    : std_logic_vector(15 downto 0);
    signal H_ADDR_A_s   : std_logic_vector(9 downto 0);
    signal H_ADDR_B_s   : std_logic_vector(9 downto 0);
    signal H_enable_B_s : std_ulogic;

begin
    -- the main program

    -- Y memory signals
	 Y_ADDR_A_s <= "00"&Y_i;
    Y_ADDR_B_s <= "0"&adress_i(8 downto 0);
    Y_enable_B_s <=adress_i(9) and valid_i;

    -- RAMB16_S18_S18: Spartan-3 1k x 16 + 2 Parity bits Dual-Port RAM
    RAMB16_Y_inst : RAMB16_S18_S18
    generic map (
      INIT_A => X"00000", --  Value of output RAM registers at startup
      INIT_B => X"00000", --  Value of output RAM registers at startup
		SRVAL_A => X"00000", --  Ouput value upon SSR assertion
      SRVAL_B => X"00000", --  Ouput value upon SSR assertion
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
		-- PORT A: Threshold
      DOA   => Y_thres_s,     -- 16-bit Data Output
      DOPA  => open,          -- 2-bit parity Output
      ADDRA => Y_ADDR_A_s,    -- 10-bit Address Input
      CLKA  => clk_i,         -- Clock
      DIA   => X"0000",       -- 16-bit Data Input
      DIPA  => "00",          -- 2-bit parity Input
      ENA   => '1',           -- RAM Enable Input
      SSRA  => '0',           -- Synchronous Set/Reset Input
      WEA   => '0',           -- Write Enable Input
		
		-- PORT B: modification
      DOB   => open,          -- 16-bit Data Output
      DOPB  => open,          -- 2-bit parity Output
      ADDRB => Y_ADDR_B_s,    -- 10-bit Address Input
      CLKB  => clk_i,         -- Clock
      DIB   => value_i,       -- 16-bit Data Input
      DIPB  => "00",          -- 2-bit parity Input
      ENB   => Y_enable_B_s,  -- RAM Enable Input
      SSRB  => '0',           -- Synchronous Set/Reset Input
      WEB   => '1'            -- Write Enable Input
    ); 
	 
	 
   -- H memory signals
	 H_ADDR_A_s <= "00"&H_i;
    H_ADDR_B_s <= "0"&adress_i(8 downto 0);
    H_enable_B_s <=not(adress_i(9)) and valid_i;

    -- RAMB16_S18_S18: Spartan-3 1k x 16 + 2 Parity bits Dual-Port RAM
    RAMB16_H_inst : RAMB16_S18_S18
    generic map (
      INIT_A => X"00000", --  Value of output RAM registers at startup
      INIT_B => X"00000", --  Value of output RAM registers at startup
		SRVAL_A => X"00000", --  Ouput value upon SSR assertion
      SRVAL_B => X"00000", --  Ouput value upon SSR assertion
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
		-- PORT A: Threshold
      DOA   => H_thres_s,     -- 16-bit Data Output
      DOPA  => open,          -- 2-bit parity Output
      ADDRA => H_ADDR_A_s,    -- 10-bit Address Input
      CLKA  => clk_i,         -- Clock
      DIA   => X"0000",       -- 16-bit Data Input
      DIPA  => "00",          -- 2-bit parity Input
      ENA   => '1',           -- RAM Enable Input
      SSRA  => '0',           -- Synchronous Set/Reset Input
      WEA   => '0',           -- Write Enable Input
		
		-- PORT B: modification
      DOB   => open,          -- 16-bit Data Output
      DOPB  => open,          -- 2-bit parity Output
      ADDRB => H_ADDR_B_s,    -- 10-bit Address Input
      CLKB  => clk_i,         -- Clock
      DIB   => value_i,       -- 16-bit Data Input
      DIPB  => "00",          -- 2-bit parity Input
      ENB   => H_enable_B_s,  -- RAM Enable Input
      SSRB  => '0',           -- Synchronous Set/Reset Input
      WEB   => '1'            -- Write Enable Input
    ); 
	 
    -- output = true => H_thres_s && Y_thres_s
    latch_out_p : process
	 begin
        wait until rising_edge(clk_i);
		  result_o <= H_thres_s and Y_thres_s;
    end process latch_out_p;
	 
end threshold_1; 
